<svg width="394" height="220" viewBox="0 0 394 220" fill="none" xmlns="http://www.w3.org/2000/svg">
<g filter="url(#filter0_d_1_858)">
<rect width="382.777" height="205.231" rx="102.615" fill="white" shape-rendering="crispEdges"/>
<rect x="7" y="7" width="368.777" height="191.231" rx="95.6153" stroke="#3A3A3A" stroke-width="14" shape-rendering="crispEdges"/>
<path d="M160.019 98.3069C161.96 103.277 162.348 107.975 161.184 112.401C160.019 116.75 157.806 120.594 154.544 123.933C151.283 127.194 147.4 129.835 142.896 131.854C138.47 133.795 134.004 134.921 129.5 135.232C126.006 135.62 122.55 135.193 119.134 133.95C115.717 132.63 112.844 130.572 110.514 127.777C108.262 124.904 107.214 121.642 107.369 117.992C107.679 111.314 107.874 101.84 107.951 89.5707C108.107 77.3012 108.223 69.5746 108.301 66.3907C108.378 64.9153 108.728 63.5175 109.349 62.1974C110.048 60.8773 110.902 59.7901 111.912 58.9359C112.999 58.004 114.241 57.2275 115.639 56.6062C117.115 55.9073 118.512 55.3638 119.832 54.9755C121.23 54.5096 122.628 54.1601 124.026 53.9271C127.287 53.4612 130.471 53.3447 133.577 53.5777C136.761 53.8107 139.712 54.5096 142.43 55.6744C145.148 56.7615 147.633 58.1205 149.885 59.7513C152.215 61.3044 154.078 63.2457 155.476 65.5754C156.951 67.905 157.961 70.3511 158.505 72.9137C159.126 75.3987 159.126 78.1943 158.505 81.3005C157.883 84.329 156.641 87.3964 154.777 90.5026C154.777 90.4249 155.127 90.852 155.825 91.7839C156.524 92.6381 157.301 93.7252 158.155 95.0454C159.087 96.3655 159.708 97.4527 160.019 98.3069ZM128.685 74.8939C128.607 76.2917 128.569 79.9803 128.569 85.9597C133.461 83.8631 136.567 81.2616 137.887 78.1554C138.586 76.7577 138.159 75.787 136.606 75.2434C135.053 74.6998 133.344 74.4668 131.481 74.5445C129.617 74.6221 128.685 74.7386 128.685 74.8939ZM140.916 107.392C141.304 106.383 141.032 105.839 140.1 105.762C139.479 105.762 137.654 106.072 134.626 106.694C131.675 107.237 129.462 107.742 127.986 108.208V114.964C129.617 114.653 130.937 114.343 131.947 114.032C132.956 113.721 134.121 113.294 135.441 112.751C136.761 112.129 137.887 111.392 138.819 110.537C139.751 109.606 140.45 108.557 140.916 107.392ZM221.901 66.5072C222.056 68.9145 222.056 71.7877 221.901 75.1269C221.901 76.2141 221.823 78.6602 221.668 82.4653C221.513 86.2704 221.357 88.9883 221.202 90.619C221.124 92.2498 220.93 94.7736 220.62 98.1904C220.309 101.607 219.882 104.325 219.338 106.344C218.795 108.363 218.096 110.732 217.242 113.45C216.387 116.09 215.3 118.497 213.98 120.671C212.66 122.846 211.107 124.865 209.321 126.729C205.438 131 200.818 133.64 195.459 134.649C190.179 135.581 185.131 134.843 180.317 132.436C175.502 129.951 171.775 126.107 169.134 120.904C167.038 116.556 165.485 111.896 164.475 106.927C163.543 101.957 163.194 96.8702 163.427 91.6674C163.66 86.3869 164.126 81.4946 164.825 76.9906C165.524 72.4866 166.494 67.5167 167.737 62.0809C168.203 59.5959 169.29 57.6157 170.998 56.1403C172.784 54.5872 174.726 53.733 176.822 53.5777C178.919 53.4224 180.938 53.6554 182.879 54.2766C184.898 54.8202 186.49 56.0238 187.655 57.8875C188.898 59.7513 189.364 61.9644 189.053 64.527C188.898 65.6919 188.509 68.4098 187.888 72.6808C187.267 76.9518 186.84 79.9803 186.607 81.7664C186.451 83.5524 186.257 86.1539 186.024 89.5707C185.791 92.9099 185.753 95.9772 185.908 98.7728C186.063 101.491 186.413 104.209 186.956 106.927C187.189 108.169 187.655 109.411 188.354 110.654C189.131 111.819 189.985 112.595 190.917 112.984C191.926 113.372 192.974 112.789 194.062 111.236C195.615 108.518 196.585 106.15 196.974 104.131C198.527 95.4336 199.769 82.6982 200.701 65.9248C201.012 62.8963 202.254 60.5666 204.429 58.9359C206.603 57.3051 208.933 56.5286 211.417 56.6062C213.98 56.6839 216.31 57.6157 218.406 59.4018C220.581 61.1102 221.746 63.4787 221.901 66.5072ZM243.038 63.4787C243.271 64.2552 243.698 65.8083 244.319 68.138C245.018 70.39 245.6 72.2537 246.066 73.7291C246.532 75.1269 247.115 76.7188 247.814 78.5049C248.513 80.2133 249.173 81.5334 249.794 82.4653C254.375 69.1863 256.86 62.0032 257.249 60.9161C258.724 56.5674 261.481 54.0048 265.519 53.2283C269.091 52.4517 272.197 53.3836 274.837 56.0238C277.555 58.5864 278.526 61.6538 277.75 65.2259C277.672 65.6918 276.235 70.0793 273.44 78.3884C270.722 86.6198 268.198 95.1618 265.868 104.014C263.616 112.867 262.49 119.623 262.49 124.282C262.413 126.845 261.675 129.097 260.277 131.038C258.957 132.902 257.171 134.106 254.919 134.649C251.968 135.348 249.522 135.309 247.581 134.533C245.639 133.679 244.242 132.553 243.387 131.155C242.533 129.679 241.99 127.544 241.757 124.748C241.601 121.953 241.601 119.701 241.757 117.992C241.912 116.206 242.145 113.799 242.455 110.77C242.455 110.537 242.455 110.382 242.455 110.305C242.533 110.149 242.572 109.994 242.572 109.839C242.572 109.606 242.611 109.411 242.688 109.256C242.844 107.625 242.378 106.422 241.291 105.645C238.65 103.626 236.282 101.219 234.185 98.4233C232.089 95.5501 230.341 92.4051 228.944 88.9883C227.546 85.5715 226.381 82.3488 225.449 79.3203C224.517 76.2141 223.663 72.7584 222.886 68.9534C222.498 66.5461 222.809 64.3717 223.818 62.4303C224.828 60.489 226.226 59.0912 228.012 58.237C229.875 57.3051 231.778 56.7615 233.719 56.6062C235.738 56.4509 237.602 56.9945 239.31 58.237C241.096 59.4795 242.339 61.2267 243.038 63.4787Z" fill="#3A3A3A"/>
</g>
<defs>
<filter id="filter0_d_1_858" x="0" y="0" width="393.871" height="219.097" filterUnits="userSpaceOnUse" color-interpolation-filters="sRGB">
<feFlood flood-opacity="0" result="BackgroundImageFix"/>
<feColorMatrix in="SourceAlpha" type="matrix" values="0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 127 0" result="hardAlpha"/>
<feOffset dx="11.0935" dy="13.8669"/>
<feComposite in2="hardAlpha" operator="out"/>
<feColorMatrix type="matrix" values="0 0 0 0 0.666667 0 0 0 0 0.290196 0 0 0 0 0.219608 0 0 0 1 0"/>
<feBlend mode="normal" in2="BackgroundImageFix" result="effect1_dropShadow_1_858"/>
<feBlend mode="normal" in="SourceGraphic" in2="effect1_dropShadow_1_858" result="shape"/>
</filter>
</defs>
</svg>
